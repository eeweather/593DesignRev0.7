module tb;

top_hdl DUT();

initial begin
   DUT.m_if.system_reset();
end

endmodule
