/*  ECE593 Project 2023wi
*   Victoria Van Gaasbeck <vvan@pdx.edu>
*   Julia Filipchuk <bfilipc2@pdx.edu>
*   Emily Weatherford <ew22@pdx.edu>
*   Daniel Keller <dk27@pdx.edu>
*
*   ALU sequence for generating ALU sequences 
*/

class sequence_alu extends uvm_sequence #(item_base);
	`uvm_object_utils(sequence_alu)

    item_base tx;

	function new(string name="sequence_alu");
		super.new(name);
	endfunction

	agent_config agent_cfg;

	task init_start(input uvm_sequencer #(item_base) sqr, input agent_config agent_cfg);
		this.agent_cfg = agent_cfg;
		this.start(sqr);
	endtask: init_start

	//generate a sequence of 10 ALU transactions
	task body();
		
		repeat (10) begin
			tx = item_alu::type_id::create("tx");
			start_item(tx);
			if(!tx.randomize()) `uvm_fatal(get_type_name(), "tx.randomize failed")
			finish_item(tx);
		end		
	
	endtask: body

endclass: sequence_alu